--==============================================================================
-- Company        : Synchrotron SOLEIL
-- Project        : PandABox FPGA
-- Design name    : sfp_udp_complete
-- Module name    : sfp_udp_complete_component_pkg.vhd
-- Purpose        : package of components declarations
-- Author         : created automatically
-- Synthesizable  : YES
-- Language       : VHDL-93
--------------------------------------------------------------------------------
-- Copyright (c) 2021 Synchrotron SOLEIL - L'Orme des Merisiers Saint-Aubin
-- BP 48 91192 Gif-sur-Yvette Cedex  - https://www.synchrotron-soleil.fr
--------------------------------------------------------------------------------
-- IMPORTANT  : THIS FILE IS AUTOMATICALLY GENERATED FROM ENTITIES LIST
--              DO NOT MODIFY IT.
--==============================================================================


--==============================================================================
-- Libraries Declaration
--==============================================================================
library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

library work;
  use work.axi_types.all;
  use work.ipv4_types.all;
  use work.arp_types.all;
  use work.top_defines.all;


--==============================================================================
-- Package Declaration
--==============================================================================
package sfp_udp_complete_component_pkg is

  component udp_complete_ping_nomac
    generic (
      CLOCK_FREQ              : integer := 125000000  ; -- freq of data_in_clk -- needed to timout cntr
      ARP_TIMEOUT             : integer := 60         ; -- ARP response timeout (s)
      ARP_MAX_PKT_TMO         : integer := 5          ; -- # wrong nwk pkts received before set error
      MAX_ARP_ENTRIES         : integer := 255        ; -- max entries in the ARP store
      --
      NB_TX_CHANNELS          : integer := 2            -- number of ip_tx channels (2 to C_MAX_CHANNELS)
    );
    port (
      -- System signals (in)
      rx_clk                  : in  std_logic;
      tx_clk                  : in  std_logic;
      reset                   : in  std_logic;
      our_ip_address          : in  std_logic_vector(31 downto 0);
      our_mac_address         : in  std_logic_vector(47 downto 0);
      control                 : in  udp_control_type;
      -- Status signals (out)
      arp_pkt_count           : out std_logic_vector(7 downto 0);   -- count of arp pkts received
      ip_pkt_count            : out std_logic_vector(7 downto 0);   -- number of IP pkts received for us
      icmp_pkt_count          : out std_logic_vector(7 downto 0);   -- number of ICMP pkts received for us
      -- UDP TX signals (in)
      udp_tx_start            : in  std_logic;                      -- indicates req to tx UDP
      udp_txi                 : in  udp_tx_type;                    -- UDP tx cxns
      udp_tx_result           : out std_logic_vector(1 downto 0);   -- tx status (changes during transmission)
      udp_tx_data_out_ready   : out std_logic;                      -- indicates udp_tx is ready to take data
      -- UDP RX signals (out)
      udp_rx_start            : out std_logic;                      -- indicates receipt of udp header
      udp_rxo                 : out udp_rx_type;
      -- IP RX signals (out)
      ip_rx_start             : out std_logic;        -- DEBUG
      ip_rx_hdr               : out ipv4_rx_header_type;
      ip_rx_data              : out axi_in_type;     -- DEBUG
      -- MAC Receiver (in)
      mac_rx_tdata            : in  std_logic_vector(7 downto 0);   -- data byte received
      mac_rx_tvalid           : in  std_logic;                      -- indicates tdata is valid
      mac_rx_tready           : out std_logic;                      -- tells mac that we are ready to take data
      mac_rx_tlast            : in  std_logic;                      -- indicates last byte of the trame
      -- MAC Transmitter (out)
      mac_tx_tdata            : out std_logic_vector(7 downto 0);   -- data byte to tx
      mac_tx_tvalid           : out std_logic;                      -- tdata is valid
      mac_tx_tready           : in  std_logic;                      -- mac is ready to accept data
      mac_tx_tfirst           : out std_logic;                      -- indicates first byte of frame
      mac_tx_tlast            : out std_logic                       -- indicates last byte of frame
    );
  end component;

  component tri_mode_ethernet_mac_0_fifo_block
     port(
        gtx_clk                    : in  std_logic;
        -- asynchronous reset
        glbl_rstn                  : in  std_logic;
        rx_axi_rstn                : in  std_logic;
        tx_axi_rstn                : in  std_logic;
        -- Reference clock for IDELAYCTRL's
        --refclk                     : in  std_logic;
        -- Receiver Statistics Interface
        -----------------------------------------
        rx_mac_aclk                : out std_logic;
        rx_reset                   : out std_logic;
        rx_statistics_vector       : out std_logic_vector(27 downto 0);
        rx_statistics_valid        : out std_logic;
        -- Receiver (AXI-S) Interface
        ------------------------------------------
        rx_fifo_clock              : in  std_logic;
        rx_fifo_resetn             : in  std_logic;
        rx_axis_fifo_tdata         : out std_logic_vector(7 downto 0);
        rx_axis_fifo_tvalid        : out std_logic;
        rx_axis_fifo_tready        : in  std_logic;
        rx_axis_fifo_tlast         : out std_logic;
        -- Transmitter Statistics Interface
        --------------------------------------------
        tx_mac_aclk                : out std_logic;
        tx_reset                   : out std_logic;
        tx_ifg_delay               : in  std_logic_vector(7 downto 0);
        tx_statistics_vector       : out std_logic_vector(31 downto 0);
        tx_statistics_valid        : out std_logic;
        -- Transmitter (AXI-S) Interface
        ---------------------------------------------
        tx_fifo_clock              : in  std_logic;
        tx_fifo_resetn             : in  std_logic;
        tx_axis_fifo_tdata         : in  std_logic_vector(7 downto 0);
        tx_axis_fifo_tvalid        : in  std_logic;
        tx_axis_fifo_tready        : out std_logic;
        tx_axis_fifo_tlast         : in  std_logic;
        tx_fifo_overflow           : out std_logic;
        tx_fifo_status             : out std_logic_vector(3 downto 0);
        -- MAC Control Interface
        --------------------------
        pause_req                  : in  std_logic;
        pause_val                  : in  std_logic_vector(15 downto 0);
        -- GMII Interface
        -------------------
        gmii_txd                  : out std_logic_vector(7 downto 0);
        gmii_tx_en                : out std_logic;
        gmii_tx_er                : out std_logic;
        gmii_tx_clk               : out std_logic;
        gmii_rxd                  : in  std_logic_vector(7 downto 0);
        gmii_rx_dv                : in  std_logic;
        gmii_rx_er                : in  std_logic;
        gmii_rx_clk               : in  std_logic;
        -- Configuration Vector
        -------------------------
        rx_configuration_vector   : in  std_logic_vector(79 downto 0);
        tx_configuration_vector   : in  std_logic_vector(79 downto 0)
     );
  end component;

  component gig_ethernet_pcs_pma_0_example_design
        port(
        -- Tranceiver Interface
        -----------------------
        gtrefclk             : in std_logic;
        gtrefclk_bufg        : in std_logic;
        txoutclk             : out std_logic;
        rxoutclk             : out std_logic;
        resetdone            : out std_logic;                    -- The GT transceiver has completed its reset cycle
        cplllock             : out std_logic;
        mmcm_reset           : out std_logic;
        mmcm_locked          : in std_logic;                     -- Locked indication from MMCM
        userclk              : in std_logic;
        userclk2             : in std_logic;
        rxuserclk              : in std_logic;
        rxuserclk2             : in std_logic;
        independent_clock_bufg : in std_logic;
        pma_reset            : in std_logic;                     -- transceiver PMA reset signal
        txp                  : out std_logic;                    -- Differential +ve of serial transmission from PMA to PMD.
        txn                  : out std_logic;                    -- Differential -ve of serial transmission from PMA to PMD.
        rxp                  : in std_logic;                     -- Differential +ve for serial reception from PMD to PMA.
        rxn                  : in std_logic;                     -- Differential -ve for serial reception from PMD to PMA.
        -- GMII Interface (client MAC <=> PCS)
        --------------------------------------
        gmii_tx_clk          : in std_logic;                     -- Transmit clock from client MAC.
        gmii_rx_clk          : out std_logic;                    -- Receive clock to client MAC.
        gmii_txd             : in std_logic_vector(7 downto 0);  -- Transmit data from client MAC.
        gmii_tx_en           : in std_logic;                     -- Transmit control signal from client MAC.
        gmii_tx_er           : in std_logic;                     -- Transmit control signal from client MAC.
        gmii_rxd             : out std_logic_vector(7 downto 0); -- Received Data to client MAC.
        gmii_rx_dv           : out std_logic;                    -- Received control signal to client MAC.
        gmii_rx_er           : out std_logic;                    -- Received control signal to client MAC.
        -- Management: Alternative to MDIO Interface
        --------------------------------------------
        configuration_vector : in std_logic_vector(4 downto 0);  -- Alternative to MDIO interface.
        -- General IO's
        ---------------
        status_vector        : out std_logic_vector(15 downto 0); -- Core status.
        reset                : in std_logic;                      -- Asynchronous reset for entire core.
        signal_detect        : in std_logic;                      -- Input from PMD to indicate presence of optical input.
        gt0_qplloutclk       : in std_logic;
        gt0_qplloutrefclk    : in std_logic
        );
  end component;

  component gig_ethernet_pcs_pma_0_clocking
     port (
        gtrefclk                : in  std_logic;                -- Reference clock for MGT: 125MHz, very high quality.
        txoutclk                : in  std_logic;                -- txoutclk from GT transceiver.
        rxoutclk                : in  std_logic;                -- rxoutclk from GT transceiver.
        mmcm_reset              : in  std_logic;                -- MMCM Reset
        gtrefclk_bufg           : out std_logic;                -- gtrefclk routed through a BUFG for driving logic.
        mmcm_locked             : out std_logic;                -- MMCM locked
        userclk                 : out std_logic;                -- for GT PMA reference clock
        userclk2                : out std_logic;                 -- 125MHz clock for core reference clock.
        rxuserclk               : out std_logic;                -- for GT PMA reference clock
        rxuserclk2              : out std_logic                 -- 125MHz clock for core reference clock.
     );
  end component;

  component gig_ethernet_pcs_pma_0_resets
     port (
      reset                    : in  std_logic;                -- Asynchronous reset for entire core.
      independent_clock_bufg   : in  std_logic;                -- System clock
      pma_reset                : out std_logic                 -- Synchronous transcevier PMA reset
     );
  end component;

  component gig_ethernet_pcs_pma_0_gt_common
  generic
  (
      -- Simulation attributes
      WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE"        -- Set to "true" to speed up sim reset
  );
  port
  (
      GTREFCLK0_IN : in std_logic;
      QPLLLOCK_OUT : out std_logic;
      QPLLLOCKDETCLK_IN : in std_logic;
      QPLLOUTCLK_OUT : out std_logic;
      QPLLOUTREFCLK_OUT : out std_logic;
      QPLLREFCLKLOST_OUT : out std_logic;
      QPLLRESET_IN : in std_logic
  );
  end component;

end sfp_udp_complete_component_pkg;

--==============================================================================
-- Package Body
--==============================================================================
package body sfp_udp_complete_component_pkg is

end package body sfp_udp_complete_component_pkg;
--==============================================================================
-- Package End
--==============================================================================
