--==============================================================================
-- Company        : Synchrotron SOLEIL
-- Project        : PandABox FPGA
-- Design name    : sfp_udpontrig
-- Module name    : udp_layer_component_pkg.vhd
-- Purpose        : package of components declarations for UDP layer
-- Author         : created automatically
-- Synthesizable  : YES
-- Language       : VHDL-93
--------------------------------------------------------------------------------
-- Copyright (c) 2021 Synchrotron SOLEIL - L'Orme des Merisiers Saint-Aubin
-- BP 48 91192 Gif-sur-Yvette Cedex  - https://www.synchrotron-soleil.fr
--------------------------------------------------------------------------------
-- IMPORTANT  : THIS FILE IS AUTOMATICALLY GENERATED FROM ENTITIES LIST
--              DO NOT MODIFY IT.
--==============================================================================


--==============================================================================
-- Libraries Declaration
--==============================================================================
library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

library work;
  use work.axi_types.all;
  use work.arp_types.all;
  use work.ipv4_types.all;
  use work.ipv4_channels_types.all;


--==============================================================================
-- Package Declaration
--==============================================================================
package udp_layer_component_pkg is

  component ip_complete_nomac
    generic (
      use_arpv2             : boolean := FALSE      ;   -- use ARP with multipule entries.
                                                        -- for single entry, set to FALSE
      no_default_gateway    : boolean := FALSE      ;   -- set to FALSE if communicating with devices accessed
                                                        -- through a "default gateway or router"
      CLOCK_FREQ            : integer := 125000000  ;   -- freq of data_in_clk -- needed to timout cntr
      ARP_TIMEOUT           : integer := 60         ;   -- ARP response timeout (s)
      ARP_MAX_PKT_TMO       : integer := 5          ;   -- # wrong nwk pkts received before set error
      MAX_ARP_ENTRIES       : integer := 255            -- max entries in the ARP store
      );
    port (
      -- IP Layer TX signals (in)
      ip_tx_start           : in  std_logic;
      ip_tx                 : in  ipv4_tx_type;                   -- IP tx cxns
      ip_tx_result          : out std_logic_vector (1 downto 0);  -- tx status (changes during transmission)
      ip_tx_data_out_ready  : out std_logic;                      -- indicates IP TX is ready to take data
      -- IP layer RX signals (out)
      ip_rx_start           : out std_logic;                      -- indicates receipt of ip frame.
      ip_rx                 : out ipv4_rx_type;
      -- system signals
      rx_clk                : in  std_logic;
      tx_clk                : in  std_logic;
      reset                 : in  std_logic;
      our_ip_address        : in  std_logic_vector (31 downto 0);
      our_mac_address       : in  std_logic_vector (47 downto 0);
      control               : in  ip_control_type;
      -- status signals
      arp_pkt_count         : out std_logic_vector(7 downto 0);   -- count of arp pkts received
      ip_pkt_count          : out std_logic_vector(7 downto 0);   -- number of IP pkts received for us
      -- MAC Transmitter
      mac_tx_tdata          : out std_logic_vector(7 downto 0);   -- data byte to tx
      mac_tx_tvalid         : out std_logic;                      -- tdata is valid
      mac_tx_tready         : in  std_logic;                      -- mac is ready to accept data
      mac_tx_tfirst         : out std_logic;                      -- indicates first byte of frame
      mac_tx_tlast          : out std_logic;                      -- indicates last byte of frame
      -- MAC Receiver
      mac_rx_tdata          : in  std_logic_vector(7 downto 0);   -- data byte received
      mac_rx_tvalid         : in  std_logic;                      -- indicates tdata is valid
      mac_rx_tready         : out std_logic;                      -- tells mac that we are ready to take data
      mac_rx_tlast          : in  std_logic                       -- indicates last byte of the trame
      );
  end component;

  component ip_tx_arbitrator
    generic (
      NB_CHANNELS               : integer := 2       -- nb of ip_tx channels (2 to C_MAX_CHANNELS)
    );
    port (
      -- System signals (in)
      clk                     : in  std_logic;                      -- asynchronous clock
      reset                   : in  std_logic;                      -- synchronous active high reset input
      -- IP layer TX input channels (in)
      ip_tx_start_bus         : in  ip_tx_start_array(0 to NB_CHANNELS-1);
      ip_tx_bus               : in  ip_tx_bus_array(0 to NB_CHANNELS-1);
      ip_tx_result_bus        : out ip_tx_result_array(0 to NB_CHANNELS-1);
      ip_tx_dout_ready_bus    : out ip_tx_dout_ready_array(0 to NB_CHANNELS-1);
     -- IP layer TX signals (out)
      ip_tx_start             : out  std_logic;
      ip_tx                   : out ipv4_tx_type;                   -- IP tx cxns
      ip_tx_result            : in  std_logic_vector(1 downto 0);   -- tx status (changes during transmission)
      ip_tx_data_out_ready    : in  std_logic                       -- indicates IP TX is ready to take data
    );
  end component;

  component udp_ping
    generic (
      -- Limit the amount of logic cells used to store ICMP optional data (synthesis only)
      -- Windows ping issues 32 bytes of ICMP data by default
      -- Linux   ping issues 64 bytes of ICMP data by default (8 bytes of header & 56 bytes of optional data)
      -- Theoritical max ping size with non fragmented IPv4 frames is 1472 bytes, ie 1500 - 20 (Ipv4 header) -8 (icmp header)
      MAX_PING_SIZE         : natural := 1024  -- 256                    -- Maximum pkt size. Larger echo requests will be ignored. (max 1472)
    );
    port (
      -- System signals (in)
      clk                   : in  std_logic;                      -- asynchronous clock
      reset                 : in  std_logic;                      -- synchronous active high reset input
      -- IP layer RX signals (in)
      ip_rx_start           : in  std_logic;                      -- indicates receipt of ip frame
      ip_rx                 : in  ipv4_rx_type;                   -- IP rx cxns
      -- status signals (out)
      icmp_pkt_count        : out std_logic_vector(7 downto 0);   -- number of ICMP pkts received for us
      icmp_pkt_err          : out std_logic;                      -- indicate an errored ICMP pkt (type <> x"0800" or pkt greater than 1472 bytes)
      icmp_pkt_err_count    : out std_logic_vector(7 downto 0);   -- number of errored ICMP pkts received for us
      -- IP layer TX signals (out)
      ip_tx_start           : out  std_logic;
      ip_tx                 : out ipv4_tx_type;                   -- IP tx cxns
      ip_tx_result          : in  std_logic_vector(1 downto 0);   -- tx status (changes during transmission)
      ip_tx_data_out_ready  : in  std_logic                       -- indicates IP TX is ready to take data
      );
  end component;

  component udp_tx
    port (
      -- system signals (in)
      clk                     : in  std_logic;                      -- same clock used to clock mac data and ip data
      reset                   : in  std_logic;
      -- UDP Layer signals (in)
      udp_tx_start            : in  std_logic;                      -- indicates req to tx UDP
      udp_txi                 : in  udp_tx_type;                    -- UDP tx cxns
      udp_tx_result           : out std_logic_vector (1 downto 0);  -- tx status (changes during transmission)
      udp_tx_data_out_ready   : out std_logic;                      -- indicates udp_tx is ready to take data
      -- IP layer TX signals (out)
      ip_tx_start             : out std_logic;
      ip_tx                   : out ipv4_tx_type;                   -- IP tx cxns
      ip_tx_result            : in  std_logic_vector (1 downto 0);  -- tx status (changes during transmission)
      ip_tx_data_out_ready    : in  std_logic                       -- indicates IP TX is ready to take data
      );
  end component;

  component udp_rx
    port (
      -- system signals
      clk             : in  std_logic;
      reset           : in  std_logic;
      -- IP layer RX signals (in)
      ip_rx_start     : in  std_logic;       -- indicates receipt of ip header
      ip_rx           : in  ipv4_rx_type;
      -- UDP Layer signals (out)
      udp_rx_start    : out std_logic;       -- indicates receipt of udp header
      udp_rxo         : out udp_rx_type
      );
  end component;

end udp_layer_component_pkg;

--==============================================================================
-- Package Body
--==============================================================================
package body udp_layer_component_pkg is

end package body udp_layer_component_pkg;
--==============================================================================
-- Package End
--==============================================================================
