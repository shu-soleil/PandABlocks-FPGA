--==============================================================================
-- Company        : Synchrotron SOLEIL
-- Project        : PandABox FPGA
-- Design name    : sfp_udpontrig
-- Module name    : ipv4_component_pkg.vhd
-- Purpose        : package of components declarations
-- Author         : created automatically
-- Synthesizable  : YES
-- Language       : VHDL-93
--------------------------------------------------------------------------------
-- Copyright (c) 2021 Synchrotron SOLEIL - L'Orme des Merisiers Saint-Aubin
-- BP 48 91192 Gif-sur-Yvette Cedex  - https://www.synchrotron-soleil.fr
--------------------------------------------------------------------------------
-- IMPORTANT  : THIS FILE IS AUTOMATICALLY GENERATED FROM ENTITIES LIST
--              DO NOT MODIFY IT.
--==============================================================================


--==============================================================================
-- Libraries Declaration
--==============================================================================
library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

library work;
  use work.axi_types.all;
  use work.ipv4_types.all;
  use work.arp_types.all;


--==============================================================================
-- Package Declaration
--==============================================================================
package ipv4_component_pkg is

  component ipv4_tx
    port (
      -- IP Layer signals
      ip_tx_start           : in  std_logic;
      ip_tx                 : in  ipv4_tx_type;                   -- IP tx cxns
      ip_tx_result          : out std_logic_vector(1 downto 0);  -- tx status (changes during transmission)
      ip_tx_data_out_ready  : out std_logic;                      -- indicates IP TX is ready to take data
      -- system signals
      clk                   : in  std_logic;                      -- same clock used to clock mac data and ip data
      reset                 : in  std_logic;
      our_ip_address        : in  std_logic_vector(31 downto 0);
      our_mac_address       : in  std_logic_vector(47 downto 0);
      -- ARP lookup signals
      arp_req_req           : out arp_req_req_type;
      arp_req_rslt          : in  arp_req_rslt_type;
      -- MAC layer TX signals
      mac_tx_req            : out std_logic;                      -- indicates that ip wants access to channel (stays up for as long as tx)
      mac_tx_granted        : in  std_logic;                      -- indicates that access to channel has been granted
      mac_data_out_ready    : in  std_logic;                      -- indicates system ready to consume data
      mac_data_out_valid    : out std_logic;                      -- indicates data out is valid
      mac_data_out_first    : out std_logic;                      -- with data out valid indicates the first byte of a frame
      mac_data_out_last     : out std_logic;                      -- with data out valid indicates the last byte of a frame
      mac_data_out          : out std_logic_vector(7 downto 0)    -- ethernet frame (from dst mac addr through to last byte of frame)
      );
  end component;

  component ipv4_rx
    port (
      -- IP Layer signals
      ip_rx             : out ipv4_rx_type;
      ip_rx_start       : out std_logic;                      -- indicates receipt of ip frame.
      -- system signals
      clk               : in  std_logic;                      -- same clock used to clock mac data and ip data
      reset             : in  std_logic;
      our_ip_address    : in  std_logic_vector(31 downto 0);
      rx_pkt_count      : out std_logic_vector( 7 downto 0);  -- number of IP pkts received for us
      -- MAC layer RX signals
      mac_data_in       : in  std_logic_vector( 7 downto 0);  -- ethernet frame (from dst mac addr through to last byte of frame)
      mac_data_in_valid : in  std_logic;                      -- indicates data_in valid on clock
      mac_data_in_last  : in  std_logic                       -- indicates last data in frame
      );
  end component;

end ipv4_component_pkg;

--==============================================================================
-- Package Body
--==============================================================================
package body ipv4_component_pkg is

end package body ipv4_component_pkg;
--==============================================================================
-- Package End
--==============================================================================
